module RegConst(
		output reg [4:0] Const29,
		output reg [4:0] Const30,
		output reg [4:0] Const31
	);
	always @(*) begin
		Const29 = 5'd29;
		Const30 = 5'd30;
		Const31 = 5'd31;
	end
endmodule
