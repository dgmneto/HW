module ULAConst(
		output reg [31:0] Const4
	);
	always @(*) 
		Const4 = 32'd4;
endmodule
